library ieee;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity VGA_image_generator is
PORT(
clock: in STD_LOGIC;
VGA_input: in STD_LOGIC_VECTOR(6 downto 0);
color_Red: out STD_LOGIC_VECTOR(3 downto 0);
color_Green: out STD_LOGIC_VECTOR(3 downto 0);
color_Blue: out STD_LOGIC_VECTOR(3 downto 0);
H_S: out STD_LOGIC;
V_S: out STD_LOGIC
);
end VGA_image_generator;


Architecture Behavioral of VGA_image_generator IS
type letter_A_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_A : letter_A_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000011000000000000000",
"00000000000000011000000000000000",
"00000000000000111100000000000000",
"00000000000000100110000000000000",
"00000000000000100110000000000000",
"00000000000001100110000000000000",
"00000000000001100010000000000000",
"00000000000001000011000000000000",
"00000000000011000001100000000000",
"00000000000110000001100000000000",
"00000000000110000001100000000000",
"00000000000110000001110000000000",
"00000000000111111111110000000000",
"00000000001100000000011000000000",
"00000000001100000000011000000000",
"00000000011000000000011000000000",
"00000000011000000000011100000000",
"00000000011000000000001100000000",
"00000000110000000000000110000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

type letter_B_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_B : letter_B_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000111111111111000000000",
"00000000000110000001111000000000",
"00000000000110000000001100000000",
"00000000000110000000001100000000",
"00000000000110000000001100000000",
"00000000000110000000001100000000",
"00000000000110000000011000000000",
"00000000000110000001100000000000",
"00000000000111111111110000000000",
"00000000000110000000011100000000",
"00000000000110000000000110000000",
"00000000000110000000000111000000",
"00000000000110000000000111000000",
"00000000000110000000000111000000",
"00000000000110000000000111000000",
"00000000000110000000000111000000",
"00000000000110000000000110000000",
"00000000000111111111111100000000",
"00000000000111111111110000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

type letter_C_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_C : letter_C_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000001111111100000000000",
"00000000000111111111111100000000",
"00000000011110000000011110000000",
"00000000111000000000000111000000",
"00000001110000000000000011100000",
"00000011110000000000000011100000",
"00000011100000000000000011000000",
"00000011000000000000000000000000",
"00000111000000000000000000000000",
"00000111000000000000000000000000",
"00000111000000000000000000000000",
"00000111000000000000000000000000",
"00000111000000000000000000000000",
"00000111000000000000000000000000",
"00000111000000000000000000000000",
"00000011100000000000000000000000",
"00000011100000000000000011100000",
"00000011110000000000000011100000",
"00000001110000000000000011100000",
"00000000111100000000001111000000",
"00000000001111000001111100000000",
"00000000001111111111111100000000",
"00000000000001111111100000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

type letter_D_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_D : letter_D_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000010000000000000000000000",
"00000000111110000000000000000000",
"00000000111111000000000000000000",
"00000000111111111000000000000000",
"00000000110000111110000000000000",
"00000000110000011111000000000000",
"00000000110000000111100000000000",
"00000000110000000001111000000000",
"00000000110000000000111000000000",
"00000000110000000000011100000000",
"00000000110000000000000110000000",
"00000000110000000000000111000000",
"00000000110000000000000111000000",
"00000000110000000000000011000000",
"00000000110000000000000011000000",
"00000000110000000000000011000000",
"00000000110000000000000011000000",
"00000000110000000000000011000000",
"00000000110000000000000011000000",
"00000000110000000000000111000000",
"00000000110000000000000111000000",
"00000000110000000000001110000000",
"00000000110000000000011100000000",
"00000000111000000000111000000000",
"00000000111111111111110000000000",
"00000000001111111111000000000000",
"00000000000011111100000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

type letter_E_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_E : letter_E_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000011111111111110000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011111111111110000000000",
"00000000011111111111110000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011000000000000000000000",
"00000000011111111111111000000000",
"00000000011111111111111000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

type letter_F_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_F : letter_F_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000001110000000000",
"00000000000111111111111000000000",
"00000000000111111111111000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000111111111100000000000",
"00000000000111111111100000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000110000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

type letter_G_array is array(0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
constant letter_G : letter_G_array :=("00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000001111100000000000",
"00000000000011110000011111000000",
"00000000000110000000000011100000",
"00000000001100000000000000100000",
"00000000001000000000000000000000",
"00000000011000000000000000000000",
"00000000111000000000000000000000",
"00000000110000000000000000000000",
"00000000110000000000000000000000",
"00000001110000000000000000000000",
"00000001110000000000000000000000",
"00000001110000000000000000000000",
"00000001110000000000111111100000",
"00000001110000000000000001100000",
"00000000110000000000000001100000",
"00000000110000000000000001100000",
"00000000111000000000000001100000",
"00000000011000000000000001100000",
"00000000001000000000000001100000",
"00000000001100000000000001100000",
"00000000000111000000000011100000",
"00000000000011110000001111000000",
"00000000000001111111111100000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

-----1280x1024 @ 60 Hz pixel clock 
signal position_h: INTEGER RANGE 0 TO 800:=0;
signal position_v: INTEGER RANGE 0 TO 525:=0;
begin

process(clock)
begin
IF(Clock'EVENT AND Clock='1')then
     
IF(VGA_input(0)='0')then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_A(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'1');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
	END IF;
    END IF;
    
if (VGA_input(1)='0') then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_B(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'1');
color_Green <= (others =>'1');
color_Blue <=(others =>'0');
end if;
end if;

if (VGA_input(2)='0') then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_C(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'0');
color_Green <= (others =>'1');
color_Blue <=(others =>'0');
end if;
end if;

if (VGA_input(3)='0') then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_D(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'0');
color_Green <= (others =>'1');
color_Blue <=(others =>'1');
end if;
end if;

if (VGA_input(4)='0') then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_E(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'1');
end if;
end if;

if (VGA_input(5)='0') then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_F(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'1');
color_Green <= (others =>'0');
color_Blue <=(others =>'1');
end if;
end if;

if (VGA_input(6)='0') then
elsif ((position_h>=144 and position_h<784) and( position_v>=33 and position_v<513)) then			
if letter_G(position_v-33)(639-(position_h-144)) = '0' then
color_Red <= (others =>'0');
color_Green <= (others =>'0');
color_Blue <=(others =>'0');
else
color_Red <= (others =>'1');
color_Green <= (others =>'1');
color_Blue <=(others =>'1');
end if;
end if;
  		
		if(position_h<800)then
		position_h<=position_h+1;
		else
		position_h<=0;
		if(position_v<525)then
	    position_v<=position_v+1;
		else
	    position_v<=0;  
		end if;  		     
		end if;
   if((position_h>0 AND position_h<160) OR (position_v>0 AND position_v<45))then
	color_Red <=(others=>'0');
	color_Green <=(others=>'0');
	color_Blue <=(others=>'0');
	end if;
   if(position_h>16 AND position_h<112)then
	   H_S<='0';
	else
	   H_S<='1';
	end if;
   if(position_v>0 AND position_v<12)then
	   V_S<='0';
	else
	   V_S<='1';
	end if;
 end if;
 end process;
 end Behavioral;